// nios_system.v

// Generated using ACDS version 15.1 189

`timescale 1 ps / 1 ps
module nios_system (
		output wire [10:0] address_export,    //    address.export
		output wire        char_read_export,  //  char_read.export
		input  wire        char_recv_export,  //  char_recv.export
		input  wire        char_sent_export,  //  char_sent.export
		output wire        chipreset_export,  //  chipreset.export
		input  wire        clk_clk,           //        clk.clk
		inout  wire [7:0]  data_export,       //       data.export
		input  wire [7:0]  data_in_export,    //    data_in.export
		output wire [7:0]  data_out_export,   //   data_out.export
		output wire [7:0]  leds_export,       //       leds.export
		output wire        load_export,       //       load.export
		output wire        notouten_export,   //   notouten.export
		output wire        readnwrite_export, // readnwrite.export
		input  wire        reset_reset_n,     //      reset.reset_n
		output wire        trans_en_export,   //   trans_en.export
		output wire [7:0]  yourboard0_export, // yourboard0.export
		output wire [7:0]  yourboard1_export, // yourboard1.export
		output wire [7:0]  yourboard2_export, // yourboard2.export
		output wire [7:0]  yourboard3_export, // yourboard3.export
		output wire [7:0]  yourboard4_export, // yourboard4.export
		output wire [7:0]  yourboard5_export, // yourboard5.export
		output wire [7:0]  yourboard6_export, // yourboard6.export
		output wire [7:0]  yourboard7_export, // yourboard7.export
		output wire [7:0]  yourshots0_export, // yourshots0.export
		output wire [7:0]  yourshots1_export, // yourshots1.export
		output wire [7:0]  yourshots2_export, // yourshots2.export
		output wire [7:0]  yourshots3_export, // yourshots3.export
		output wire [7:0]  yourshots4_export, // yourshots4.export
		output wire [7:0]  yourshots5_export, // yourshots5.export
		output wire [7:0]  yourshots6_export, // yourshots6.export
		output wire [7:0]  yourshots7_export  // yourshots7.export
	);

	wire  [31:0] nios2_processor_data_master_readdata;                            // mm_interconnect_0:nios2_processor_data_master_readdata -> nios2_processor:d_readdata
	wire         nios2_processor_data_master_waitrequest;                         // mm_interconnect_0:nios2_processor_data_master_waitrequest -> nios2_processor:d_waitrequest
	wire         nios2_processor_data_master_debugaccess;                         // nios2_processor:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_processor_data_master_debugaccess
	wire  [17:0] nios2_processor_data_master_address;                             // nios2_processor:d_address -> mm_interconnect_0:nios2_processor_data_master_address
	wire   [3:0] nios2_processor_data_master_byteenable;                          // nios2_processor:d_byteenable -> mm_interconnect_0:nios2_processor_data_master_byteenable
	wire         nios2_processor_data_master_read;                                // nios2_processor:d_read -> mm_interconnect_0:nios2_processor_data_master_read
	wire         nios2_processor_data_master_write;                               // nios2_processor:d_write -> mm_interconnect_0:nios2_processor_data_master_write
	wire  [31:0] nios2_processor_data_master_writedata;                           // nios2_processor:d_writedata -> mm_interconnect_0:nios2_processor_data_master_writedata
	wire  [31:0] nios2_processor_instruction_master_readdata;                     // mm_interconnect_0:nios2_processor_instruction_master_readdata -> nios2_processor:i_readdata
	wire         nios2_processor_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_processor_instruction_master_waitrequest -> nios2_processor:i_waitrequest
	wire  [17:0] nios2_processor_instruction_master_address;                      // nios2_processor:i_address -> mm_interconnect_0:nios2_processor_instruction_master_address
	wire         nios2_processor_instruction_master_read;                         // nios2_processor:i_read -> mm_interconnect_0:nios2_processor_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;          // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;       // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_processor_jtag_debug_module_readdata;    // nios2_processor:jtag_debug_module_readdata -> mm_interconnect_0:nios2_processor_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_waitrequest; // nios2_processor:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_processor_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_processor_jtag_debug_module_debugaccess -> nios2_processor:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_processor_jtag_debug_module_address;     // mm_interconnect_0:nios2_processor_jtag_debug_module_address -> nios2_processor:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_read;        // mm_interconnect_0:nios2_processor_jtag_debug_module_read -> nios2_processor:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_processor_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_processor_jtag_debug_module_byteenable -> nios2_processor:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_write;       // mm_interconnect_0:nios2_processor_jtag_debug_module_write -> nios2_processor:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_processor_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_processor_jtag_debug_module_writedata -> nios2_processor:jtag_debug_module_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                   // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                     // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory_s1_address;                      // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                   // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                        // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                    // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                        // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_leds_s1_chipselect;                            // mm_interconnect_0:LEDs_s1_chipselect -> LEDs:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                              // LEDs:readdata -> mm_interconnect_0:LEDs_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                               // mm_interconnect_0:LEDs_s1_address -> LEDs:address
	wire         mm_interconnect_0_leds_s1_write;                                 // mm_interconnect_0:LEDs_s1_write -> LEDs:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                             // mm_interconnect_0:LEDs_s1_writedata -> LEDs:writedata
	wire         mm_interconnect_0_data_out_s1_chipselect;                        // mm_interconnect_0:data_out_s1_chipselect -> data_out:chipselect
	wire  [31:0] mm_interconnect_0_data_out_s1_readdata;                          // data_out:readdata -> mm_interconnect_0:data_out_s1_readdata
	wire   [1:0] mm_interconnect_0_data_out_s1_address;                           // mm_interconnect_0:data_out_s1_address -> data_out:address
	wire         mm_interconnect_0_data_out_s1_write;                             // mm_interconnect_0:data_out_s1_write -> data_out:write_n
	wire  [31:0] mm_interconnect_0_data_out_s1_writedata;                         // mm_interconnect_0:data_out_s1_writedata -> data_out:writedata
	wire         mm_interconnect_0_trans_en_s1_chipselect;                        // mm_interconnect_0:trans_en_s1_chipselect -> trans_en:chipselect
	wire  [31:0] mm_interconnect_0_trans_en_s1_readdata;                          // trans_en:readdata -> mm_interconnect_0:trans_en_s1_readdata
	wire   [1:0] mm_interconnect_0_trans_en_s1_address;                           // mm_interconnect_0:trans_en_s1_address -> trans_en:address
	wire         mm_interconnect_0_trans_en_s1_write;                             // mm_interconnect_0:trans_en_s1_write -> trans_en:write_n
	wire  [31:0] mm_interconnect_0_trans_en_s1_writedata;                         // mm_interconnect_0:trans_en_s1_writedata -> trans_en:writedata
	wire  [31:0] mm_interconnect_0_char_sent_s1_readdata;                         // char_sent:readdata -> mm_interconnect_0:char_sent_s1_readdata
	wire   [1:0] mm_interconnect_0_char_sent_s1_address;                          // mm_interconnect_0:char_sent_s1_address -> char_sent:address
	wire         mm_interconnect_0_load_s1_chipselect;                            // mm_interconnect_0:load_s1_chipselect -> load:chipselect
	wire  [31:0] mm_interconnect_0_load_s1_readdata;                              // load:readdata -> mm_interconnect_0:load_s1_readdata
	wire   [1:0] mm_interconnect_0_load_s1_address;                               // mm_interconnect_0:load_s1_address -> load:address
	wire         mm_interconnect_0_load_s1_write;                                 // mm_interconnect_0:load_s1_write -> load:write_n
	wire  [31:0] mm_interconnect_0_load_s1_writedata;                             // mm_interconnect_0:load_s1_writedata -> load:writedata
	wire  [31:0] mm_interconnect_0_data_in_s1_readdata;                           // data_in:readdata -> mm_interconnect_0:data_in_s1_readdata
	wire   [1:0] mm_interconnect_0_data_in_s1_address;                            // mm_interconnect_0:data_in_s1_address -> data_in:address
	wire  [31:0] mm_interconnect_0_char_recv_s1_readdata;                         // char_recv:readdata -> mm_interconnect_0:char_recv_s1_readdata
	wire   [1:0] mm_interconnect_0_char_recv_s1_address;                          // mm_interconnect_0:char_recv_s1_address -> char_recv:address
	wire         mm_interconnect_0_char_read_s1_chipselect;                       // mm_interconnect_0:char_read_s1_chipselect -> char_read:chipselect
	wire  [31:0] mm_interconnect_0_char_read_s1_readdata;                         // char_read:readdata -> mm_interconnect_0:char_read_s1_readdata
	wire   [1:0] mm_interconnect_0_char_read_s1_address;                          // mm_interconnect_0:char_read_s1_address -> char_read:address
	wire         mm_interconnect_0_char_read_s1_write;                            // mm_interconnect_0:char_read_s1_write -> char_read:write_n
	wire  [31:0] mm_interconnect_0_char_read_s1_writedata;                        // mm_interconnect_0:char_read_s1_writedata -> char_read:writedata
	wire         mm_interconnect_0_notouten_s1_chipselect;                        // mm_interconnect_0:notOutEn_s1_chipselect -> notOutEn:chipselect
	wire  [31:0] mm_interconnect_0_notouten_s1_readdata;                          // notOutEn:readdata -> mm_interconnect_0:notOutEn_s1_readdata
	wire   [1:0] mm_interconnect_0_notouten_s1_address;                           // mm_interconnect_0:notOutEn_s1_address -> notOutEn:address
	wire         mm_interconnect_0_notouten_s1_write;                             // mm_interconnect_0:notOutEn_s1_write -> notOutEn:write_n
	wire  [31:0] mm_interconnect_0_notouten_s1_writedata;                         // mm_interconnect_0:notOutEn_s1_writedata -> notOutEn:writedata
	wire         mm_interconnect_0_readnwrite_s1_chipselect;                      // mm_interconnect_0:readnWrite_s1_chipselect -> readnWrite:chipselect
	wire  [31:0] mm_interconnect_0_readnwrite_s1_readdata;                        // readnWrite:readdata -> mm_interconnect_0:readnWrite_s1_readdata
	wire   [1:0] mm_interconnect_0_readnwrite_s1_address;                         // mm_interconnect_0:readnWrite_s1_address -> readnWrite:address
	wire         mm_interconnect_0_readnwrite_s1_write;                           // mm_interconnect_0:readnWrite_s1_write -> readnWrite:write_n
	wire  [31:0] mm_interconnect_0_readnwrite_s1_writedata;                       // mm_interconnect_0:readnWrite_s1_writedata -> readnWrite:writedata
	wire         mm_interconnect_0_chipreset_s1_chipselect;                       // mm_interconnect_0:chipReset_s1_chipselect -> chipReset:chipselect
	wire  [31:0] mm_interconnect_0_chipreset_s1_readdata;                         // chipReset:readdata -> mm_interconnect_0:chipReset_s1_readdata
	wire   [1:0] mm_interconnect_0_chipreset_s1_address;                          // mm_interconnect_0:chipReset_s1_address -> chipReset:address
	wire         mm_interconnect_0_chipreset_s1_write;                            // mm_interconnect_0:chipReset_s1_write -> chipReset:write_n
	wire  [31:0] mm_interconnect_0_chipreset_s1_writedata;                        // mm_interconnect_0:chipReset_s1_writedata -> chipReset:writedata
	wire         mm_interconnect_0_address_s1_chipselect;                         // mm_interconnect_0:address_s1_chipselect -> address:chipselect
	wire  [31:0] mm_interconnect_0_address_s1_readdata;                           // address:readdata -> mm_interconnect_0:address_s1_readdata
	wire   [1:0] mm_interconnect_0_address_s1_address;                            // mm_interconnect_0:address_s1_address -> address:address
	wire         mm_interconnect_0_address_s1_write;                              // mm_interconnect_0:address_s1_write -> address:write_n
	wire  [31:0] mm_interconnect_0_address_s1_writedata;                          // mm_interconnect_0:address_s1_writedata -> address:writedata
	wire         mm_interconnect_0_data_s1_chipselect;                            // mm_interconnect_0:data_s1_chipselect -> data:chipselect
	wire  [31:0] mm_interconnect_0_data_s1_readdata;                              // data:readdata -> mm_interconnect_0:data_s1_readdata
	wire   [1:0] mm_interconnect_0_data_s1_address;                               // mm_interconnect_0:data_s1_address -> data:address
	wire         mm_interconnect_0_data_s1_write;                                 // mm_interconnect_0:data_s1_write -> data:write_n
	wire  [31:0] mm_interconnect_0_data_s1_writedata;                             // mm_interconnect_0:data_s1_writedata -> data:writedata
	wire         mm_interconnect_0_yourboard1_s1_chipselect;                      // mm_interconnect_0:yourboard1_s1_chipselect -> yourboard1:chipselect
	wire  [31:0] mm_interconnect_0_yourboard1_s1_readdata;                        // yourboard1:readdata -> mm_interconnect_0:yourboard1_s1_readdata
	wire   [1:0] mm_interconnect_0_yourboard1_s1_address;                         // mm_interconnect_0:yourboard1_s1_address -> yourboard1:address
	wire         mm_interconnect_0_yourboard1_s1_write;                           // mm_interconnect_0:yourboard1_s1_write -> yourboard1:write_n
	wire  [31:0] mm_interconnect_0_yourboard1_s1_writedata;                       // mm_interconnect_0:yourboard1_s1_writedata -> yourboard1:writedata
	wire         mm_interconnect_0_yourboard2_s1_chipselect;                      // mm_interconnect_0:yourboard2_s1_chipselect -> yourboard2:chipselect
	wire  [31:0] mm_interconnect_0_yourboard2_s1_readdata;                        // yourboard2:readdata -> mm_interconnect_0:yourboard2_s1_readdata
	wire   [1:0] mm_interconnect_0_yourboard2_s1_address;                         // mm_interconnect_0:yourboard2_s1_address -> yourboard2:address
	wire         mm_interconnect_0_yourboard2_s1_write;                           // mm_interconnect_0:yourboard2_s1_write -> yourboard2:write_n
	wire  [31:0] mm_interconnect_0_yourboard2_s1_writedata;                       // mm_interconnect_0:yourboard2_s1_writedata -> yourboard2:writedata
	wire         mm_interconnect_0_yourboard3_s1_chipselect;                      // mm_interconnect_0:yourboard3_s1_chipselect -> yourboard3:chipselect
	wire  [31:0] mm_interconnect_0_yourboard3_s1_readdata;                        // yourboard3:readdata -> mm_interconnect_0:yourboard3_s1_readdata
	wire   [1:0] mm_interconnect_0_yourboard3_s1_address;                         // mm_interconnect_0:yourboard3_s1_address -> yourboard3:address
	wire         mm_interconnect_0_yourboard3_s1_write;                           // mm_interconnect_0:yourboard3_s1_write -> yourboard3:write_n
	wire  [31:0] mm_interconnect_0_yourboard3_s1_writedata;                       // mm_interconnect_0:yourboard3_s1_writedata -> yourboard3:writedata
	wire         mm_interconnect_0_yourboard4_s1_chipselect;                      // mm_interconnect_0:yourboard4_s1_chipselect -> yourboard4:chipselect
	wire  [31:0] mm_interconnect_0_yourboard4_s1_readdata;                        // yourboard4:readdata -> mm_interconnect_0:yourboard4_s1_readdata
	wire   [1:0] mm_interconnect_0_yourboard4_s1_address;                         // mm_interconnect_0:yourboard4_s1_address -> yourboard4:address
	wire         mm_interconnect_0_yourboard4_s1_write;                           // mm_interconnect_0:yourboard4_s1_write -> yourboard4:write_n
	wire  [31:0] mm_interconnect_0_yourboard4_s1_writedata;                       // mm_interconnect_0:yourboard4_s1_writedata -> yourboard4:writedata
	wire         mm_interconnect_0_yourboard6_s1_chipselect;                      // mm_interconnect_0:yourboard6_s1_chipselect -> yourboard6:chipselect
	wire  [31:0] mm_interconnect_0_yourboard6_s1_readdata;                        // yourboard6:readdata -> mm_interconnect_0:yourboard6_s1_readdata
	wire   [1:0] mm_interconnect_0_yourboard6_s1_address;                         // mm_interconnect_0:yourboard6_s1_address -> yourboard6:address
	wire         mm_interconnect_0_yourboard6_s1_write;                           // mm_interconnect_0:yourboard6_s1_write -> yourboard6:write_n
	wire  [31:0] mm_interconnect_0_yourboard6_s1_writedata;                       // mm_interconnect_0:yourboard6_s1_writedata -> yourboard6:writedata
	wire         mm_interconnect_0_yourboard7_s1_chipselect;                      // mm_interconnect_0:yourboard7_s1_chipselect -> yourboard7:chipselect
	wire  [31:0] mm_interconnect_0_yourboard7_s1_readdata;                        // yourboard7:readdata -> mm_interconnect_0:yourboard7_s1_readdata
	wire   [1:0] mm_interconnect_0_yourboard7_s1_address;                         // mm_interconnect_0:yourboard7_s1_address -> yourboard7:address
	wire         mm_interconnect_0_yourboard7_s1_write;                           // mm_interconnect_0:yourboard7_s1_write -> yourboard7:write_n
	wire  [31:0] mm_interconnect_0_yourboard7_s1_writedata;                       // mm_interconnect_0:yourboard7_s1_writedata -> yourboard7:writedata
	wire         mm_interconnect_0_yourboard0_s1_chipselect;                      // mm_interconnect_0:yourboard0_s1_chipselect -> yourboard0:chipselect
	wire  [31:0] mm_interconnect_0_yourboard0_s1_readdata;                        // yourboard0:readdata -> mm_interconnect_0:yourboard0_s1_readdata
	wire   [1:0] mm_interconnect_0_yourboard0_s1_address;                         // mm_interconnect_0:yourboard0_s1_address -> yourboard0:address
	wire         mm_interconnect_0_yourboard0_s1_write;                           // mm_interconnect_0:yourboard0_s1_write -> yourboard0:write_n
	wire  [31:0] mm_interconnect_0_yourboard0_s1_writedata;                       // mm_interconnect_0:yourboard0_s1_writedata -> yourboard0:writedata
	wire         mm_interconnect_0_yourboard5_s1_chipselect;                      // mm_interconnect_0:yourboard5_s1_chipselect -> yourboard5:chipselect
	wire  [31:0] mm_interconnect_0_yourboard5_s1_readdata;                        // yourboard5:readdata -> mm_interconnect_0:yourboard5_s1_readdata
	wire   [1:0] mm_interconnect_0_yourboard5_s1_address;                         // mm_interconnect_0:yourboard5_s1_address -> yourboard5:address
	wire         mm_interconnect_0_yourboard5_s1_write;                           // mm_interconnect_0:yourboard5_s1_write -> yourboard5:write_n
	wire  [31:0] mm_interconnect_0_yourboard5_s1_writedata;                       // mm_interconnect_0:yourboard5_s1_writedata -> yourboard5:writedata
	wire         mm_interconnect_0_yourshots0_s1_chipselect;                      // mm_interconnect_0:yourshots0_s1_chipselect -> yourshots0:chipselect
	wire  [31:0] mm_interconnect_0_yourshots0_s1_readdata;                        // yourshots0:readdata -> mm_interconnect_0:yourshots0_s1_readdata
	wire   [1:0] mm_interconnect_0_yourshots0_s1_address;                         // mm_interconnect_0:yourshots0_s1_address -> yourshots0:address
	wire         mm_interconnect_0_yourshots0_s1_write;                           // mm_interconnect_0:yourshots0_s1_write -> yourshots0:write_n
	wire  [31:0] mm_interconnect_0_yourshots0_s1_writedata;                       // mm_interconnect_0:yourshots0_s1_writedata -> yourshots0:writedata
	wire         mm_interconnect_0_yourshots1_s1_chipselect;                      // mm_interconnect_0:yourshots1_s1_chipselect -> yourshots1:chipselect
	wire  [31:0] mm_interconnect_0_yourshots1_s1_readdata;                        // yourshots1:readdata -> mm_interconnect_0:yourshots1_s1_readdata
	wire   [1:0] mm_interconnect_0_yourshots1_s1_address;                         // mm_interconnect_0:yourshots1_s1_address -> yourshots1:address
	wire         mm_interconnect_0_yourshots1_s1_write;                           // mm_interconnect_0:yourshots1_s1_write -> yourshots1:write_n
	wire  [31:0] mm_interconnect_0_yourshots1_s1_writedata;                       // mm_interconnect_0:yourshots1_s1_writedata -> yourshots1:writedata
	wire         mm_interconnect_0_yourshots2_s1_chipselect;                      // mm_interconnect_0:yourshots2_s1_chipselect -> yourshots2:chipselect
	wire  [31:0] mm_interconnect_0_yourshots2_s1_readdata;                        // yourshots2:readdata -> mm_interconnect_0:yourshots2_s1_readdata
	wire   [1:0] mm_interconnect_0_yourshots2_s1_address;                         // mm_interconnect_0:yourshots2_s1_address -> yourshots2:address
	wire         mm_interconnect_0_yourshots2_s1_write;                           // mm_interconnect_0:yourshots2_s1_write -> yourshots2:write_n
	wire  [31:0] mm_interconnect_0_yourshots2_s1_writedata;                       // mm_interconnect_0:yourshots2_s1_writedata -> yourshots2:writedata
	wire         mm_interconnect_0_yourshots3_s1_chipselect;                      // mm_interconnect_0:yourshots3_s1_chipselect -> yourshots3:chipselect
	wire  [31:0] mm_interconnect_0_yourshots3_s1_readdata;                        // yourshots3:readdata -> mm_interconnect_0:yourshots3_s1_readdata
	wire   [1:0] mm_interconnect_0_yourshots3_s1_address;                         // mm_interconnect_0:yourshots3_s1_address -> yourshots3:address
	wire         mm_interconnect_0_yourshots3_s1_write;                           // mm_interconnect_0:yourshots3_s1_write -> yourshots3:write_n
	wire  [31:0] mm_interconnect_0_yourshots3_s1_writedata;                       // mm_interconnect_0:yourshots3_s1_writedata -> yourshots3:writedata
	wire         mm_interconnect_0_yourshots4_s1_chipselect;                      // mm_interconnect_0:yourshots4_s1_chipselect -> yourshots4:chipselect
	wire  [31:0] mm_interconnect_0_yourshots4_s1_readdata;                        // yourshots4:readdata -> mm_interconnect_0:yourshots4_s1_readdata
	wire   [1:0] mm_interconnect_0_yourshots4_s1_address;                         // mm_interconnect_0:yourshots4_s1_address -> yourshots4:address
	wire         mm_interconnect_0_yourshots4_s1_write;                           // mm_interconnect_0:yourshots4_s1_write -> yourshots4:write_n
	wire  [31:0] mm_interconnect_0_yourshots4_s1_writedata;                       // mm_interconnect_0:yourshots4_s1_writedata -> yourshots4:writedata
	wire         mm_interconnect_0_yourshots5_s1_chipselect;                      // mm_interconnect_0:yourshots5_s1_chipselect -> yourshots5:chipselect
	wire  [31:0] mm_interconnect_0_yourshots5_s1_readdata;                        // yourshots5:readdata -> mm_interconnect_0:yourshots5_s1_readdata
	wire   [1:0] mm_interconnect_0_yourshots5_s1_address;                         // mm_interconnect_0:yourshots5_s1_address -> yourshots5:address
	wire         mm_interconnect_0_yourshots5_s1_write;                           // mm_interconnect_0:yourshots5_s1_write -> yourshots5:write_n
	wire  [31:0] mm_interconnect_0_yourshots5_s1_writedata;                       // mm_interconnect_0:yourshots5_s1_writedata -> yourshots5:writedata
	wire         mm_interconnect_0_yourshots6_s1_chipselect;                      // mm_interconnect_0:yourshots6_s1_chipselect -> yourshots6:chipselect
	wire  [31:0] mm_interconnect_0_yourshots6_s1_readdata;                        // yourshots6:readdata -> mm_interconnect_0:yourshots6_s1_readdata
	wire   [1:0] mm_interconnect_0_yourshots6_s1_address;                         // mm_interconnect_0:yourshots6_s1_address -> yourshots6:address
	wire         mm_interconnect_0_yourshots6_s1_write;                           // mm_interconnect_0:yourshots6_s1_write -> yourshots6:write_n
	wire  [31:0] mm_interconnect_0_yourshots6_s1_writedata;                       // mm_interconnect_0:yourshots6_s1_writedata -> yourshots6:writedata
	wire         mm_interconnect_0_yourshots7_s1_chipselect;                      // mm_interconnect_0:yourshots7_s1_chipselect -> yourshots7:chipselect
	wire  [31:0] mm_interconnect_0_yourshots7_s1_readdata;                        // yourshots7:readdata -> mm_interconnect_0:yourshots7_s1_readdata
	wire   [1:0] mm_interconnect_0_yourshots7_s1_address;                         // mm_interconnect_0:yourshots7_s1_address -> yourshots7:address
	wire         mm_interconnect_0_yourshots7_s1_write;                           // mm_interconnect_0:yourshots7_s1_write -> yourshots7:write_n
	wire  [31:0] mm_interconnect_0_yourshots7_s1_writedata;                       // mm_interconnect_0:yourshots7_s1_writedata -> yourshots7:writedata
	wire         irq_mapper_receiver0_irq;                                        // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_processor_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_processor:d_irq
	wire         rst_controller_reset_out_reset;                                  // rst_controller:reset_out -> [LEDs:reset_n, address:reset_n, chipReset:reset_n, data:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_processor_reset_n_reset_bridge_in_reset_reset, nios2_processor:reset_n, notOutEn:reset_n, onchip_memory:reset, readnWrite:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                              // rst_controller:reset_req -> [nios2_processor:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         nios2_processor_jtag_debug_module_reset_reset;                   // nios2_processor:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                              // rst_controller_001:reset_out -> [char_read:reset_n, char_recv:reset_n, char_sent:reset_n, data_in:reset_n, data_out:reset_n, load:reset_n, mm_interconnect_0:data_out_reset_reset_bridge_in_reset_reset, trans_en:reset_n, yourboard0:reset_n, yourboard1:reset_n, yourboard2:reset_n, yourboard3:reset_n, yourboard4:reset_n, yourboard5:reset_n, yourboard6:reset_n, yourboard7:reset_n, yourshots0:reset_n, yourshots1:reset_n, yourshots2:reset_n, yourshots3:reset_n, yourshots4:reset_n, yourshots5:reset_n, yourshots6:reset_n, yourshots7:reset_n]

	nios_system_LEDs leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	nios_system_address address (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_address_s1_readdata),   //                    .readdata
		.out_port   (address_export)                           // external_connection.export
	);

	nios_system_char_read char_read (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_char_read_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_char_read_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_char_read_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_char_read_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_char_read_s1_readdata),   //                    .readdata
		.out_port   (char_read_export)                           // external_connection.export
	);

	nios_system_char_recv char_recv (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_char_recv_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_char_recv_s1_readdata), //                    .readdata
		.in_port  (char_recv_export)                         // external_connection.export
	);

	nios_system_char_recv char_sent (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_char_sent_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_char_sent_s1_readdata), //                    .readdata
		.in_port  (char_sent_export)                         // external_connection.export
	);

	nios_system_char_read chipreset (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_chipreset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chipreset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chipreset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chipreset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chipreset_s1_readdata),   //                    .readdata
		.out_port   (chipreset_export)                           // external_connection.export
	);

	nios_system_data data (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data_s1_readdata),   //                    .readdata
		.bidir_port (data_export)                           // external_connection.export
	);

	nios_system_data_in data_in (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_data_in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_data_in_s1_readdata), //                    .readdata
		.in_port  (data_in_export)                         // external_connection.export
	);

	nios_system_LEDs data_out (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_data_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data_out_s1_readdata),   //                    .readdata
		.out_port   (data_out_export)                           // external_connection.export
	);

	nios_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	nios_system_char_read load (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_load_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_load_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_load_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_load_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_load_s1_readdata),   //                    .readdata
		.out_port   (load_export)                           // external_connection.export
	);

	nios_system_nios2_processor nios2_processor (
		.clk                                   (clk_clk),                                                         //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                              //                          .reset_req
		.d_address                             (nios2_processor_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_processor_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_processor_data_master_read),                                //                          .read
		.d_readdata                            (nios2_processor_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_processor_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_processor_data_master_write),                               //                          .write
		.d_writedata                           (nios2_processor_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_processor_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_processor_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_processor_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_processor_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_processor_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_processor_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_processor_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_processor_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_processor_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_processor_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_processor_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_processor_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_processor_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_processor_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_processor_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                 // custom_instruction_master.readra
	);

	nios_system_char_read notouten (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_notouten_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_notouten_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_notouten_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_notouten_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_notouten_s1_readdata),   //                    .readdata
		.out_port   (notouten_export)                           // external_connection.export
	);

	nios_system_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	nios_system_char_read readnwrite (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_readnwrite_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_readnwrite_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_readnwrite_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_readnwrite_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_readnwrite_s1_readdata),   //                    .readdata
		.out_port   (readnwrite_export)                           // external_connection.export
	);

	nios_system_char_read trans_en (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_trans_en_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_trans_en_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_trans_en_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_trans_en_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_trans_en_s1_readdata),   //                    .readdata
		.out_port   (trans_en_export)                           // external_connection.export
	);

	nios_system_LEDs yourboard0 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourboard0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourboard0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourboard0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourboard0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourboard0_s1_readdata),   //                    .readdata
		.out_port   (yourboard0_export)                           // external_connection.export
	);

	nios_system_LEDs yourboard1 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourboard1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourboard1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourboard1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourboard1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourboard1_s1_readdata),   //                    .readdata
		.out_port   (yourboard1_export)                           // external_connection.export
	);

	nios_system_LEDs yourboard2 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourboard2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourboard2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourboard2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourboard2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourboard2_s1_readdata),   //                    .readdata
		.out_port   (yourboard2_export)                           // external_connection.export
	);

	nios_system_LEDs yourboard3 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourboard3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourboard3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourboard3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourboard3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourboard3_s1_readdata),   //                    .readdata
		.out_port   (yourboard3_export)                           // external_connection.export
	);

	nios_system_LEDs yourboard4 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourboard4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourboard4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourboard4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourboard4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourboard4_s1_readdata),   //                    .readdata
		.out_port   (yourboard4_export)                           // external_connection.export
	);

	nios_system_LEDs yourboard5 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourboard5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourboard5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourboard5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourboard5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourboard5_s1_readdata),   //                    .readdata
		.out_port   (yourboard5_export)                           // external_connection.export
	);

	nios_system_LEDs yourboard6 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourboard6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourboard6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourboard6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourboard6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourboard6_s1_readdata),   //                    .readdata
		.out_port   (yourboard6_export)                           // external_connection.export
	);

	nios_system_LEDs yourboard7 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourboard7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourboard7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourboard7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourboard7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourboard7_s1_readdata),   //                    .readdata
		.out_port   (yourboard7_export)                           // external_connection.export
	);

	nios_system_LEDs yourshots0 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourshots0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourshots0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourshots0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourshots0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourshots0_s1_readdata),   //                    .readdata
		.out_port   (yourshots0_export)                           // external_connection.export
	);

	nios_system_LEDs yourshots1 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourshots1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourshots1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourshots1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourshots1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourshots1_s1_readdata),   //                    .readdata
		.out_port   (yourshots1_export)                           // external_connection.export
	);

	nios_system_LEDs yourshots2 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourshots2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourshots2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourshots2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourshots2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourshots2_s1_readdata),   //                    .readdata
		.out_port   (yourshots2_export)                           // external_connection.export
	);

	nios_system_LEDs yourshots3 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourshots3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourshots3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourshots3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourshots3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourshots3_s1_readdata),   //                    .readdata
		.out_port   (yourshots3_export)                           // external_connection.export
	);

	nios_system_LEDs yourshots4 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourshots4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourshots4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourshots4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourshots4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourshots4_s1_readdata),   //                    .readdata
		.out_port   (yourshots4_export)                           // external_connection.export
	);

	nios_system_LEDs yourshots5 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourshots5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourshots5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourshots5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourshots5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourshots5_s1_readdata),   //                    .readdata
		.out_port   (yourshots5_export)                           // external_connection.export
	);

	nios_system_LEDs yourshots6 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourshots6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourshots6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourshots6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourshots6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourshots6_s1_readdata),   //                    .readdata
		.out_port   (yourshots6_export)                           // external_connection.export
	);

	nios_system_LEDs yourshots7 (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_yourshots7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_yourshots7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_yourshots7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_yourshots7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_yourshots7_s1_readdata),   //                    .readdata
		.out_port   (yourshots7_export)                           // external_connection.export
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                       (clk_clk),                                                         //                                     clk_0_clk.clk
		.data_out_reset_reset_bridge_in_reset_reset          (rst_controller_001_reset_out_reset),                              //          data_out_reset_reset_bridge_in_reset.reset
		.nios2_processor_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                  // nios2_processor_reset_n_reset_bridge_in_reset.reset
		.nios2_processor_data_master_address                 (nios2_processor_data_master_address),                             //                   nios2_processor_data_master.address
		.nios2_processor_data_master_waitrequest             (nios2_processor_data_master_waitrequest),                         //                                              .waitrequest
		.nios2_processor_data_master_byteenable              (nios2_processor_data_master_byteenable),                          //                                              .byteenable
		.nios2_processor_data_master_read                    (nios2_processor_data_master_read),                                //                                              .read
		.nios2_processor_data_master_readdata                (nios2_processor_data_master_readdata),                            //                                              .readdata
		.nios2_processor_data_master_write                   (nios2_processor_data_master_write),                               //                                              .write
		.nios2_processor_data_master_writedata               (nios2_processor_data_master_writedata),                           //                                              .writedata
		.nios2_processor_data_master_debugaccess             (nios2_processor_data_master_debugaccess),                         //                                              .debugaccess
		.nios2_processor_instruction_master_address          (nios2_processor_instruction_master_address),                      //            nios2_processor_instruction_master.address
		.nios2_processor_instruction_master_waitrequest      (nios2_processor_instruction_master_waitrequest),                  //                                              .waitrequest
		.nios2_processor_instruction_master_read             (nios2_processor_instruction_master_read),                         //                                              .read
		.nios2_processor_instruction_master_readdata         (nios2_processor_instruction_master_readdata),                     //                                              .readdata
		.address_s1_address                                  (mm_interconnect_0_address_s1_address),                            //                                    address_s1.address
		.address_s1_write                                    (mm_interconnect_0_address_s1_write),                              //                                              .write
		.address_s1_readdata                                 (mm_interconnect_0_address_s1_readdata),                           //                                              .readdata
		.address_s1_writedata                                (mm_interconnect_0_address_s1_writedata),                          //                                              .writedata
		.address_s1_chipselect                               (mm_interconnect_0_address_s1_chipselect),                         //                                              .chipselect
		.char_read_s1_address                                (mm_interconnect_0_char_read_s1_address),                          //                                  char_read_s1.address
		.char_read_s1_write                                  (mm_interconnect_0_char_read_s1_write),                            //                                              .write
		.char_read_s1_readdata                               (mm_interconnect_0_char_read_s1_readdata),                         //                                              .readdata
		.char_read_s1_writedata                              (mm_interconnect_0_char_read_s1_writedata),                        //                                              .writedata
		.char_read_s1_chipselect                             (mm_interconnect_0_char_read_s1_chipselect),                       //                                              .chipselect
		.char_recv_s1_address                                (mm_interconnect_0_char_recv_s1_address),                          //                                  char_recv_s1.address
		.char_recv_s1_readdata                               (mm_interconnect_0_char_recv_s1_readdata),                         //                                              .readdata
		.char_sent_s1_address                                (mm_interconnect_0_char_sent_s1_address),                          //                                  char_sent_s1.address
		.char_sent_s1_readdata                               (mm_interconnect_0_char_sent_s1_readdata),                         //                                              .readdata
		.chipReset_s1_address                                (mm_interconnect_0_chipreset_s1_address),                          //                                  chipReset_s1.address
		.chipReset_s1_write                                  (mm_interconnect_0_chipreset_s1_write),                            //                                              .write
		.chipReset_s1_readdata                               (mm_interconnect_0_chipreset_s1_readdata),                         //                                              .readdata
		.chipReset_s1_writedata                              (mm_interconnect_0_chipreset_s1_writedata),                        //                                              .writedata
		.chipReset_s1_chipselect                             (mm_interconnect_0_chipreset_s1_chipselect),                       //                                              .chipselect
		.data_s1_address                                     (mm_interconnect_0_data_s1_address),                               //                                       data_s1.address
		.data_s1_write                                       (mm_interconnect_0_data_s1_write),                                 //                                              .write
		.data_s1_readdata                                    (mm_interconnect_0_data_s1_readdata),                              //                                              .readdata
		.data_s1_writedata                                   (mm_interconnect_0_data_s1_writedata),                             //                                              .writedata
		.data_s1_chipselect                                  (mm_interconnect_0_data_s1_chipselect),                            //                                              .chipselect
		.data_in_s1_address                                  (mm_interconnect_0_data_in_s1_address),                            //                                    data_in_s1.address
		.data_in_s1_readdata                                 (mm_interconnect_0_data_in_s1_readdata),                           //                                              .readdata
		.data_out_s1_address                                 (mm_interconnect_0_data_out_s1_address),                           //                                   data_out_s1.address
		.data_out_s1_write                                   (mm_interconnect_0_data_out_s1_write),                             //                                              .write
		.data_out_s1_readdata                                (mm_interconnect_0_data_out_s1_readdata),                          //                                              .readdata
		.data_out_s1_writedata                               (mm_interconnect_0_data_out_s1_writedata),                         //                                              .writedata
		.data_out_s1_chipselect                              (mm_interconnect_0_data_out_s1_chipselect),                        //                                              .chipselect
		.jtag_uart_avalon_jtag_slave_address                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),           //                   jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),             //                                              .write
		.jtag_uart_avalon_jtag_slave_read                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),              //                                              .read
		.jtag_uart_avalon_jtag_slave_readdata                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),          //                                              .readdata
		.jtag_uart_avalon_jtag_slave_writedata               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),         //                                              .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),       //                                              .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),        //                                              .chipselect
		.LEDs_s1_address                                     (mm_interconnect_0_leds_s1_address),                               //                                       LEDs_s1.address
		.LEDs_s1_write                                       (mm_interconnect_0_leds_s1_write),                                 //                                              .write
		.LEDs_s1_readdata                                    (mm_interconnect_0_leds_s1_readdata),                              //                                              .readdata
		.LEDs_s1_writedata                                   (mm_interconnect_0_leds_s1_writedata),                             //                                              .writedata
		.LEDs_s1_chipselect                                  (mm_interconnect_0_leds_s1_chipselect),                            //                                              .chipselect
		.load_s1_address                                     (mm_interconnect_0_load_s1_address),                               //                                       load_s1.address
		.load_s1_write                                       (mm_interconnect_0_load_s1_write),                                 //                                              .write
		.load_s1_readdata                                    (mm_interconnect_0_load_s1_readdata),                              //                                              .readdata
		.load_s1_writedata                                   (mm_interconnect_0_load_s1_writedata),                             //                                              .writedata
		.load_s1_chipselect                                  (mm_interconnect_0_load_s1_chipselect),                            //                                              .chipselect
		.nios2_processor_jtag_debug_module_address           (mm_interconnect_0_nios2_processor_jtag_debug_module_address),     //             nios2_processor_jtag_debug_module.address
		.nios2_processor_jtag_debug_module_write             (mm_interconnect_0_nios2_processor_jtag_debug_module_write),       //                                              .write
		.nios2_processor_jtag_debug_module_read              (mm_interconnect_0_nios2_processor_jtag_debug_module_read),        //                                              .read
		.nios2_processor_jtag_debug_module_readdata          (mm_interconnect_0_nios2_processor_jtag_debug_module_readdata),    //                                              .readdata
		.nios2_processor_jtag_debug_module_writedata         (mm_interconnect_0_nios2_processor_jtag_debug_module_writedata),   //                                              .writedata
		.nios2_processor_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_processor_jtag_debug_module_byteenable),  //                                              .byteenable
		.nios2_processor_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_processor_jtag_debug_module_waitrequest), //                                              .waitrequest
		.nios2_processor_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_processor_jtag_debug_module_debugaccess), //                                              .debugaccess
		.notOutEn_s1_address                                 (mm_interconnect_0_notouten_s1_address),                           //                                   notOutEn_s1.address
		.notOutEn_s1_write                                   (mm_interconnect_0_notouten_s1_write),                             //                                              .write
		.notOutEn_s1_readdata                                (mm_interconnect_0_notouten_s1_readdata),                          //                                              .readdata
		.notOutEn_s1_writedata                               (mm_interconnect_0_notouten_s1_writedata),                         //                                              .writedata
		.notOutEn_s1_chipselect                              (mm_interconnect_0_notouten_s1_chipselect),                        //                                              .chipselect
		.onchip_memory_s1_address                            (mm_interconnect_0_onchip_memory_s1_address),                      //                              onchip_memory_s1.address
		.onchip_memory_s1_write                              (mm_interconnect_0_onchip_memory_s1_write),                        //                                              .write
		.onchip_memory_s1_readdata                           (mm_interconnect_0_onchip_memory_s1_readdata),                     //                                              .readdata
		.onchip_memory_s1_writedata                          (mm_interconnect_0_onchip_memory_s1_writedata),                    //                                              .writedata
		.onchip_memory_s1_byteenable                         (mm_interconnect_0_onchip_memory_s1_byteenable),                   //                                              .byteenable
		.onchip_memory_s1_chipselect                         (mm_interconnect_0_onchip_memory_s1_chipselect),                   //                                              .chipselect
		.onchip_memory_s1_clken                              (mm_interconnect_0_onchip_memory_s1_clken),                        //                                              .clken
		.readnWrite_s1_address                               (mm_interconnect_0_readnwrite_s1_address),                         //                                 readnWrite_s1.address
		.readnWrite_s1_write                                 (mm_interconnect_0_readnwrite_s1_write),                           //                                              .write
		.readnWrite_s1_readdata                              (mm_interconnect_0_readnwrite_s1_readdata),                        //                                              .readdata
		.readnWrite_s1_writedata                             (mm_interconnect_0_readnwrite_s1_writedata),                       //                                              .writedata
		.readnWrite_s1_chipselect                            (mm_interconnect_0_readnwrite_s1_chipselect),                      //                                              .chipselect
		.trans_en_s1_address                                 (mm_interconnect_0_trans_en_s1_address),                           //                                   trans_en_s1.address
		.trans_en_s1_write                                   (mm_interconnect_0_trans_en_s1_write),                             //                                              .write
		.trans_en_s1_readdata                                (mm_interconnect_0_trans_en_s1_readdata),                          //                                              .readdata
		.trans_en_s1_writedata                               (mm_interconnect_0_trans_en_s1_writedata),                         //                                              .writedata
		.trans_en_s1_chipselect                              (mm_interconnect_0_trans_en_s1_chipselect),                        //                                              .chipselect
		.yourboard0_s1_address                               (mm_interconnect_0_yourboard0_s1_address),                         //                                 yourboard0_s1.address
		.yourboard0_s1_write                                 (mm_interconnect_0_yourboard0_s1_write),                           //                                              .write
		.yourboard0_s1_readdata                              (mm_interconnect_0_yourboard0_s1_readdata),                        //                                              .readdata
		.yourboard0_s1_writedata                             (mm_interconnect_0_yourboard0_s1_writedata),                       //                                              .writedata
		.yourboard0_s1_chipselect                            (mm_interconnect_0_yourboard0_s1_chipselect),                      //                                              .chipselect
		.yourboard1_s1_address                               (mm_interconnect_0_yourboard1_s1_address),                         //                                 yourboard1_s1.address
		.yourboard1_s1_write                                 (mm_interconnect_0_yourboard1_s1_write),                           //                                              .write
		.yourboard1_s1_readdata                              (mm_interconnect_0_yourboard1_s1_readdata),                        //                                              .readdata
		.yourboard1_s1_writedata                             (mm_interconnect_0_yourboard1_s1_writedata),                       //                                              .writedata
		.yourboard1_s1_chipselect                            (mm_interconnect_0_yourboard1_s1_chipselect),                      //                                              .chipselect
		.yourboard2_s1_address                               (mm_interconnect_0_yourboard2_s1_address),                         //                                 yourboard2_s1.address
		.yourboard2_s1_write                                 (mm_interconnect_0_yourboard2_s1_write),                           //                                              .write
		.yourboard2_s1_readdata                              (mm_interconnect_0_yourboard2_s1_readdata),                        //                                              .readdata
		.yourboard2_s1_writedata                             (mm_interconnect_0_yourboard2_s1_writedata),                       //                                              .writedata
		.yourboard2_s1_chipselect                            (mm_interconnect_0_yourboard2_s1_chipselect),                      //                                              .chipselect
		.yourboard3_s1_address                               (mm_interconnect_0_yourboard3_s1_address),                         //                                 yourboard3_s1.address
		.yourboard3_s1_write                                 (mm_interconnect_0_yourboard3_s1_write),                           //                                              .write
		.yourboard3_s1_readdata                              (mm_interconnect_0_yourboard3_s1_readdata),                        //                                              .readdata
		.yourboard3_s1_writedata                             (mm_interconnect_0_yourboard3_s1_writedata),                       //                                              .writedata
		.yourboard3_s1_chipselect                            (mm_interconnect_0_yourboard3_s1_chipselect),                      //                                              .chipselect
		.yourboard4_s1_address                               (mm_interconnect_0_yourboard4_s1_address),                         //                                 yourboard4_s1.address
		.yourboard4_s1_write                                 (mm_interconnect_0_yourboard4_s1_write),                           //                                              .write
		.yourboard4_s1_readdata                              (mm_interconnect_0_yourboard4_s1_readdata),                        //                                              .readdata
		.yourboard4_s1_writedata                             (mm_interconnect_0_yourboard4_s1_writedata),                       //                                              .writedata
		.yourboard4_s1_chipselect                            (mm_interconnect_0_yourboard4_s1_chipselect),                      //                                              .chipselect
		.yourboard5_s1_address                               (mm_interconnect_0_yourboard5_s1_address),                         //                                 yourboard5_s1.address
		.yourboard5_s1_write                                 (mm_interconnect_0_yourboard5_s1_write),                           //                                              .write
		.yourboard5_s1_readdata                              (mm_interconnect_0_yourboard5_s1_readdata),                        //                                              .readdata
		.yourboard5_s1_writedata                             (mm_interconnect_0_yourboard5_s1_writedata),                       //                                              .writedata
		.yourboard5_s1_chipselect                            (mm_interconnect_0_yourboard5_s1_chipselect),                      //                                              .chipselect
		.yourboard6_s1_address                               (mm_interconnect_0_yourboard6_s1_address),                         //                                 yourboard6_s1.address
		.yourboard6_s1_write                                 (mm_interconnect_0_yourboard6_s1_write),                           //                                              .write
		.yourboard6_s1_readdata                              (mm_interconnect_0_yourboard6_s1_readdata),                        //                                              .readdata
		.yourboard6_s1_writedata                             (mm_interconnect_0_yourboard6_s1_writedata),                       //                                              .writedata
		.yourboard6_s1_chipselect                            (mm_interconnect_0_yourboard6_s1_chipselect),                      //                                              .chipselect
		.yourboard7_s1_address                               (mm_interconnect_0_yourboard7_s1_address),                         //                                 yourboard7_s1.address
		.yourboard7_s1_write                                 (mm_interconnect_0_yourboard7_s1_write),                           //                                              .write
		.yourboard7_s1_readdata                              (mm_interconnect_0_yourboard7_s1_readdata),                        //                                              .readdata
		.yourboard7_s1_writedata                             (mm_interconnect_0_yourboard7_s1_writedata),                       //                                              .writedata
		.yourboard7_s1_chipselect                            (mm_interconnect_0_yourboard7_s1_chipselect),                      //                                              .chipselect
		.yourshots0_s1_address                               (mm_interconnect_0_yourshots0_s1_address),                         //                                 yourshots0_s1.address
		.yourshots0_s1_write                                 (mm_interconnect_0_yourshots0_s1_write),                           //                                              .write
		.yourshots0_s1_readdata                              (mm_interconnect_0_yourshots0_s1_readdata),                        //                                              .readdata
		.yourshots0_s1_writedata                             (mm_interconnect_0_yourshots0_s1_writedata),                       //                                              .writedata
		.yourshots0_s1_chipselect                            (mm_interconnect_0_yourshots0_s1_chipselect),                      //                                              .chipselect
		.yourshots1_s1_address                               (mm_interconnect_0_yourshots1_s1_address),                         //                                 yourshots1_s1.address
		.yourshots1_s1_write                                 (mm_interconnect_0_yourshots1_s1_write),                           //                                              .write
		.yourshots1_s1_readdata                              (mm_interconnect_0_yourshots1_s1_readdata),                        //                                              .readdata
		.yourshots1_s1_writedata                             (mm_interconnect_0_yourshots1_s1_writedata),                       //                                              .writedata
		.yourshots1_s1_chipselect                            (mm_interconnect_0_yourshots1_s1_chipselect),                      //                                              .chipselect
		.yourshots2_s1_address                               (mm_interconnect_0_yourshots2_s1_address),                         //                                 yourshots2_s1.address
		.yourshots2_s1_write                                 (mm_interconnect_0_yourshots2_s1_write),                           //                                              .write
		.yourshots2_s1_readdata                              (mm_interconnect_0_yourshots2_s1_readdata),                        //                                              .readdata
		.yourshots2_s1_writedata                             (mm_interconnect_0_yourshots2_s1_writedata),                       //                                              .writedata
		.yourshots2_s1_chipselect                            (mm_interconnect_0_yourshots2_s1_chipselect),                      //                                              .chipselect
		.yourshots3_s1_address                               (mm_interconnect_0_yourshots3_s1_address),                         //                                 yourshots3_s1.address
		.yourshots3_s1_write                                 (mm_interconnect_0_yourshots3_s1_write),                           //                                              .write
		.yourshots3_s1_readdata                              (mm_interconnect_0_yourshots3_s1_readdata),                        //                                              .readdata
		.yourshots3_s1_writedata                             (mm_interconnect_0_yourshots3_s1_writedata),                       //                                              .writedata
		.yourshots3_s1_chipselect                            (mm_interconnect_0_yourshots3_s1_chipselect),                      //                                              .chipselect
		.yourshots4_s1_address                               (mm_interconnect_0_yourshots4_s1_address),                         //                                 yourshots4_s1.address
		.yourshots4_s1_write                                 (mm_interconnect_0_yourshots4_s1_write),                           //                                              .write
		.yourshots4_s1_readdata                              (mm_interconnect_0_yourshots4_s1_readdata),                        //                                              .readdata
		.yourshots4_s1_writedata                             (mm_interconnect_0_yourshots4_s1_writedata),                       //                                              .writedata
		.yourshots4_s1_chipselect                            (mm_interconnect_0_yourshots4_s1_chipselect),                      //                                              .chipselect
		.yourshots5_s1_address                               (mm_interconnect_0_yourshots5_s1_address),                         //                                 yourshots5_s1.address
		.yourshots5_s1_write                                 (mm_interconnect_0_yourshots5_s1_write),                           //                                              .write
		.yourshots5_s1_readdata                              (mm_interconnect_0_yourshots5_s1_readdata),                        //                                              .readdata
		.yourshots5_s1_writedata                             (mm_interconnect_0_yourshots5_s1_writedata),                       //                                              .writedata
		.yourshots5_s1_chipselect                            (mm_interconnect_0_yourshots5_s1_chipselect),                      //                                              .chipselect
		.yourshots6_s1_address                               (mm_interconnect_0_yourshots6_s1_address),                         //                                 yourshots6_s1.address
		.yourshots6_s1_write                                 (mm_interconnect_0_yourshots6_s1_write),                           //                                              .write
		.yourshots6_s1_readdata                              (mm_interconnect_0_yourshots6_s1_readdata),                        //                                              .readdata
		.yourshots6_s1_writedata                             (mm_interconnect_0_yourshots6_s1_writedata),                       //                                              .writedata
		.yourshots6_s1_chipselect                            (mm_interconnect_0_yourshots6_s1_chipselect),                      //                                              .chipselect
		.yourshots7_s1_address                               (mm_interconnect_0_yourshots7_s1_address),                         //                                 yourshots7_s1.address
		.yourshots7_s1_write                                 (mm_interconnect_0_yourshots7_s1_write),                           //                                              .write
		.yourshots7_s1_readdata                              (mm_interconnect_0_yourshots7_s1_readdata),                        //                                              .readdata
		.yourshots7_s1_writedata                             (mm_interconnect_0_yourshots7_s1_writedata),                       //                                              .writedata
		.yourshots7_s1_chipselect                            (mm_interconnect_0_yourshots7_s1_chipselect)                       //                                              .chipselect
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_processor_d_irq_irq)       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                                // reset_in0.reset
		.reset_in1      (nios2_processor_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),                // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),            //          .reset_req
		.reset_req_in0  (1'b0),                                          // (terminated)
		.reset_req_in1  (1'b0),                                          // (terminated)
		.reset_in2      (1'b0),                                          // (terminated)
		.reset_req_in2  (1'b0),                                          // (terminated)
		.reset_in3      (1'b0),                                          // (terminated)
		.reset_req_in3  (1'b0),                                          // (terminated)
		.reset_in4      (1'b0),                                          // (terminated)
		.reset_req_in4  (1'b0),                                          // (terminated)
		.reset_in5      (1'b0),                                          // (terminated)
		.reset_req_in5  (1'b0),                                          // (terminated)
		.reset_in6      (1'b0),                                          // (terminated)
		.reset_req_in6  (1'b0),                                          // (terminated)
		.reset_in7      (1'b0),                                          // (terminated)
		.reset_req_in7  (1'b0),                                          // (terminated)
		.reset_in8      (1'b0),                                          // (terminated)
		.reset_req_in8  (1'b0),                                          // (terminated)
		.reset_in9      (1'b0),                                          // (terminated)
		.reset_req_in9  (1'b0),                                          // (terminated)
		.reset_in10     (1'b0),                                          // (terminated)
		.reset_req_in10 (1'b0),                                          // (terminated)
		.reset_in11     (1'b0),                                          // (terminated)
		.reset_req_in11 (1'b0),                                          // (terminated)
		.reset_in12     (1'b0),                                          // (terminated)
		.reset_req_in12 (1'b0),                                          // (terminated)
		.reset_in13     (1'b0),                                          // (terminated)
		.reset_req_in13 (1'b0),                                          // (terminated)
		.reset_in14     (1'b0),                                          // (terminated)
		.reset_req_in14 (1'b0),                                          // (terminated)
		.reset_in15     (1'b0),                                          // (terminated)
		.reset_req_in15 (1'b0)                                           // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
