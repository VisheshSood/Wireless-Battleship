//In & out ports consist of 8 parallel wires, an input address of 12 bits chooses the address to access in the RAM,
//and the system will either read from RAM or write to RAM based on the configuration of the
//active low input signals, "not output enable" and "read not write"

//This specific RAM consists of 2048 addresses, each containing one byte of data.

module sram (data, address, notOutEn, readnWrite, chipSelect);
    inout [7:0] data;
    input [10:0] address;
    input notOutEn, readnWrite, chipSelect;
    reg [7:0] ram [2047:0];

    assign data = (~notOutEn & ~chipSelect) ? ram[address] : 8'bz;

    //Perform the write operation when read signal is strobed high
    always @(posedge readnWrite)
        //Overwrites the memory at proper address using the input signal on the data bus
        if (~chipSelect)
            ram[address] <= data;

endmodule

